library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity default is
    Port ();
end default;

architecture Behavioral of default is



begin



end Behavioral;